//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Apr 14 19:02:26 2017
// Version: v11.7 SP1 11.7.1.14
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// touch_screen
module touch_screen(
    // Inputs
    SPI_1_DI,
    // Outputs
    SPI_1_DO,
    // Inouts
    I2C_1_SCL,
    I2C_1_SDA,
    SPI_1_CLK,
    SPI_1_SS
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  SPI_1_DI;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output SPI_1_DO;
//--------------------------------------------------------------------
// Inout
//--------------------------------------------------------------------
inout  I2C_1_SCL;
inout  I2C_1_SDA;
inout  SPI_1_CLK;
inout  SPI_1_SS;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   I2C_1_SCL;
wire   I2C_1_SDA;
wire   SPI_1_CLK;
wire   SPI_1_DI;
wire   SPI_1_DO_net_0;
wire   SPI_1_SS;
wire   SPI_1_DO_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign SPI_1_DO_net_1 = SPI_1_DO_net_0;
assign SPI_1_DO       = SPI_1_DO_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------touch_screen_MSS
touch_screen_MSS touch_screen_MSS_0(
        // Inputs
        .SPI_1_DI  ( SPI_1_DI ),
        // Outputs
        .SPI_1_DO  ( SPI_1_DO_net_0 ),
        // Inouts
        .SPI_1_CLK ( SPI_1_CLK ),
        .SPI_1_SS  ( SPI_1_SS ),
        .I2C_1_SCL ( I2C_1_SCL ),
        .I2C_1_SDA ( I2C_1_SDA ) 
        );


endmodule
